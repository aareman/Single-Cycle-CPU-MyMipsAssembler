library verilog;
use verilog.vl_types.all;
entity Instruction_man_vlg_vec_tst is
end Instruction_man_vlg_vec_tst;
