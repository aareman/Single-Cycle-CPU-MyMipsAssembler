library verilog;
use verilog.vl_types.all;
entity r_typeIn_vlg_vec_tst is
end r_typeIn_vlg_vec_tst;
