library ieee; 
use ieee.std_logic_1164.all; 
use IEEE.numeric_std.all;


entity instructionFile is     
	port (address: in std_logic_vector(4 downto 0);
			outInstruction: out std_logic_vector(31 downto 0));    -- clock and reset 
end instructionFile; 
	-- purpose: Main 	architecture details for SIMPREG 
architecture arch of instructionFile is 	
	begin  	
	-- SIMPLE     
process (address)	
type NIBBLE is array (31 downto 0) of std_logic;
	type MEM is array (0 to 31) of NIBBLE;
-- an array "array of array" type
	variable MEM32X32 : MEM;
begin	

MEM32X32(0):= "00000000000000000000000000000000";
MEM32X32(1):= "01010100000000010000000000000000";
MEM32X32(2):= "01010100000000100000000000000001";
MEM32X32(3):= "01010100000000110000000000000000";
MEM32X32(4):= "01010100000000000000000000000000";
MEM32X32(5):= "00010000010000000001100000000000";
MEM32X32(6):= "00010000010000010001000000000000";
MEM32X32(7):= "00010000011000000000100000000000";
MEM32X32(8):= "10000100010000101111111111111101";
MEM32X32(9):= "01010100000001010000000000001111";
MEM32X32(10):= "01010100000001010000000000001111";
MEM32X32(11):= "01010100000001010000000000001111";
MEM32X32(12):= "01010100000001010000000000001111";
MEM32X32(13):= "01010100000001010000000000001111";
MEM32X32(14):= "01010100000001010000000000001111";
MEM32X32(15):= "01010100000001010000000000001111";
MEM32X32(16):= "01010100000001010000000000001111";
MEM32X32(17):= "01010100000001010000000000001111";
MEM32X32(18):= "01010100000001010000000000001111";
MEM32X32(19):= "01010100000001010000000000001111";
MEM32X32(20):= "01010100000001010000000000001111";
MEM32X32(21):= "01010100000001010000000000001111";
MEM32X32(22):= "01010100000001010000000000001111";
MEM32X32(23):= "01010100000001010000000000001111";
MEM32X32(24):= "01010100000001010000000000001111";
MEM32X32(25):= "01010100000001010000000000001111";
MEM32X32(26):= "01010100000001010000000000001111";
MEM32X32(27):= "01010100000001010000000000001111";
MEM32X32(28):= "01010100000001010000000000001111";
MEM32X32(29):= "01010100000001010000000000001111";
MEM32X32(30):= "01010100000001010000000000001111";
MEM32X32(31):= "01010100000001010000000000001111";

--	MEM32X32(1):= "010101" & "00000010101111111111111111"; -- li r10, -1
--	MEM32X32(2):= "010101" & "00000101000000000000000010"; -- li r20, 2
--	MEM32X32(3):= "000100" & "10100010101111000000000000"; -- add r30, r20, r10
--	MEM32X32(4):= "100010" & "10101101011111111111111101"; -- beq r20, r20, -3
--	MEM32X32(5):= "010101" & "00000010100000000000000011"; -- li r10, 3
--	
--MEM32X32(0):= "00000000000000000000000000000000";
--MEM32X32(1):= "01010100000101000000000000001010";
--MEM32X32(2):= "01010100000000000000000000000000";
--MEM32X32(3):= "01001110100101001111111111111110";
--MEM32X32(4):= "10001010100000001111111111111111";
	outInstruction <= std_logic_vector(MEM32X32(to_integer(unsigned(address))));	
end process;

end arch;

